// ============================================================================
//  文件名   : mux2.v
//  模块名   : mux2
// ----------------------------------------------------------------------------
//  功能描述 : 可参数化位宽的 2:1 多路选择器
//             ┌────────────┐            ┌────────────┐
//             │ 输入 d0[N:0]│ ----s=0-->│            │
//             │ 输入 d1[N:0]│ ----s=1-->│    y = ?   │───► 输出 y[N:0]
//             │ 选择信号 s  │           │            │
//             └────────────┘            └────────────┘
//             • 当 s=0 时输出 d0；当 s=1 时输出 d1。
// ----------------------------------------------------------------------------
//  Verilog-2001 说明
//    1. SystemVerilog 的 `logic` 全部改为省略类型（默认 wire）。           |
//    2. 参数列表结尾 **不要** 加分号：`#(parameter WIDTH = 8)`               |
//    3. 纯组合逻辑用 `assign` 连续赋值即可，无需 `always @*`。              |
// ============================================================================
module mux2 #(
  parameter WIDTH = 8  // 数据位宽，默认 8 位
) (
  input  [WIDTH-1:0] d0,  // 输入 0
  input  [WIDTH-1:0] d1,  // 输入 1
  input              s,   // 选择信号（高选 d1，低选 d0）
  output [WIDTH-1:0] y    // 输出
);

  // --------------------------------------------------------------------
  // 组合多路选择：s=0 选 d0，s=1 选 d1
  // --------------------------------------------------------------------
  assign y = s ? d1 : d0;

endmodule
