// ============================================================================
//  文件名   : imem.v
//  模块名   : imem
// ----------------------------------------------------------------------------
//  功能描述 : 指令存储器（64 × 32-bit ROM, 读延迟 0）
//             • 地址 a 以 **字节地址** 形式给出，内部取 a[31:2] 作为字索引；
//             • 仿真时用 $readmemh 从 “memfile.dat” 把机器码预加载进 ROM；
//             • 读口 rd 为 **异步组合**，地址变化立即输出指令字。
// ----------------------------------------------------------------------------
//  Verilog-2001 迁移要点
//    1) SystemVerilog 的 `logic` → Verilog 的 `wire` / `reg`
//       ─ 端口 a/rd 默认 wire；内部存储阵列 ROM 声明为 reg。
//    2) 连续赋值 `assign rd = ROM[...]` 保持异步读行为。
//    3) ANSI-style 端口写法在 IEEE-1364-2001 已被广泛支持。
// ============================================================================
(* dont_touch = "true" *) module imem (
  input         clka,  // 时钟
  input  [31:0] a_0,     // 字节地址（来自 PC）
  output [31:0] rd_0,     // 读出指令字
  input  [31:0] a_1,     // 字节地址（来自 PC）
  output [31:0] rd_1,      // 读出指令字
  input  [31:0] a_2,     // 字节地址（来自 PC）
  output [31:0] rd_2,      // 读出指令字
  input  [31:0] a_3,     // 字节地址（来自 PC）
  output [31:0] rd_3,      // 读出指令字
  input  [31:0] a_4,     // 字节地址（来自 PC）
  output [31:0] rd_4,      // 读出指令字
  input  [31:0] a_5,     // 字节地址（来自 PC）
  output [31:0] rd_5,      // 读出指令字
  input  [31:0] a_6,     // 字节地址（来自 PC）
  output [31:0] rd_6,      // 读出指令字
  input  [31:0] a_7,     // 字节地址（来自 PC）
  output [31:0] rd_7       // 读出指令
);
  // rom ROM (
  //   .clka (clka),
  //   .addra(a[31:2]),
  //   .douta(rd)
  // );
  imem_0 ROM_1 (
    .a  (a_0[31:2]),  // input wire [6 : 0] a
    .spo(rd_0)        // output wire [31 : 0] spo
  );

  imem_1 ROM_2 (
    .a  (a_1[31:2]),  // input wire [6 : 0] a
    .spo(rd_1)        // output wire [31 : 0] spo
  );

  imem_2 ROM_3 (
    .a  (a_2[31:2]),  // input wire [6 : 0] a
    .spo(rd_2)        // output wire [31 : 0] spo
  );

  imem_3 ROM_4 (
    .a  (a_3[31:2]),  // input wire [6 : 0] a
    .spo(rd_3)        // output wire [31 : 0] spo
  );

  imem_4 ROM_5 (
    .a  (a_4[31:2]),  // input wire [6 : 0] a
    .spo(rd_4)        // output wire [31 : 0] spo
  );

  imem_5 ROM_6 (
    .a  (a_5[31:2]),  // input wire [6 : 0] a
    .spo(rd_5)        // output wire [31 : 0] spo
  );

  imem_6 ROM_7 (
    .a  (a_6[31:2]),  // input wire [6 : 0] a
    .spo(rd_6)        // output wire [31 : 0] spo
  );

  imem_7 ROM_8 (
    .a  (a_7[31:2]),  // input wire [6 : 0] a
    .spo(rd_7)        // output wire [31 : 0] spo
  );
  // --------------------------------------------------------------------
  // 64 × 32-bit 只读存储器；Synth 时综合工具会将 initial 数据固化到 ROM。
  // --------------------------------------------------------------------
  // reg [31:0] ROM[0:63];

  // --------------------------------------------------------------------
  // 初始化：仿真启动时把 “memfile.dat” 中的十六进制指令加载进 ROM。
  //   • 每行写一个 32-bit 十六进制数（不带 0x），见前文示例 prog.hex。
  // --------------------------------------------------------------------
  // initial begin
  //   $readmemh("memfile.mem", ROM);
  // end

  // --------------------------------------------------------------------
  // 异步读：地址变化立即输出，对应硬件为 “组合查表”。
  // 字对齐 → 舍弃最低 2 位（字节地址 → 字地址）
  // --------------------------------------------------------------------
  // assign rd = ROM[a[31:2]];

endmodule
