// ============================================================================
//  文件名   : dmem.v
//  模块名   : dmem
// ----------------------------------------------------------------------------
//  功能描述 : **32-bit 单端口数据存储器**（写同步、读异步）  
//             • 地址选择逻辑：
//               - a值在0-15 → 读取ROM_1
//               - a值在16-47 → 读取RAM
//               - a值在48-63 → 读取verify_RAM
// ============================================================================
module dmem (
  input         clk,  // 时钟
  input         we,   // 写使能（高有效）
  input  [31:0] a,    // 地址（字节对齐，取高位[31:2] 作索引）
  input  [31:0] wd,   // 写入数据
  output [31:0] rd    // 读出数据
);

  // --------------------------------------------------------------------
  // 1) 内部存储阵列：64 × 32-bit（可通过修改深度扩展容量）
  // --------------------------------------------------------------------
  reg  [31:0] RAM                                [47:16];
  reg  [31:0] verify_RAM                         [63:48];  // 修正命名为统一大写
  wire [15:0] rom_data;  // ROM_1 输出数据
  reg  [31:0] mem_data;  // 最终选择的数据

  // // 行为级仿真初始化
  // initial begin
  //   $readmemh("FFT_input.mem", RAM);  // 每行一字（16-bit）
  // end

  // --------------------------------------------------------------------
  // 2) 存储器读取实例
  // --------------------------------------------------------------------
  dist_mem_gen_1 ROM_1 (
    .a  (a[4:1]),   // input wire [3 : 0] a
    .spo(rom_data)  // output wire [15 : 0] spo
  );

  // --------------------------------------------------------------------
  // 3) 根据地址范围选择读取源
  // --------------------------------------------------------------------
  always @(*) begin
    if (a[8:1] <= 7'd15) begin
      // 地址范围 0-15，从ROM_1读取
      mem_data = {16'b0, rom_data};
    end else if (a[8:1] >= 7'd16 && a[8:1] <= 7'd47) begin
      // 地址范围 16-47，从RAM读取
      mem_data = {16'b0, RAM[a[8:1]]};
    end else if (a[8:1] >= 7'd48 && a[8:1] <= 7'd63) begin
      // 地址范围 48-63，从verify_RAM读取
      mem_data = {16'b0, verify_RAM[a[8:1]]};
    end else begin
      // 超出范围，返回0或其他默认值
      mem_data = 32'h0000_0000;
    end
  end

  // 输出连接到选择后的数据
  assign rd = mem_data;

  // --------------------------------------------------------------------
  // 4) 同步写入（按照需要写入对应存储器）
  // --------------------------------------------------------------------
  always @(posedge clk) begin
    if (we) begin
      if (a[8:1] >= 7'd16 && a[8:1] <= 7'd47) RAM[a[8:1]] <= wd[15:0];
      else if (a[8:1] >= 7'd48 && a[8:1] <= 7'd63) verify_RAM[a[8:1]] <= wd[15:0];
      // ROM通常不可写入，此处不处理ROM写入
    end
  end

endmodule
