`timescale 1ns / 1ps
// ============================================================================
//  文件名   : tb_imem.v
//  模块名   : tb_imem (testbench for imem)
// ----------------------------------------------------------------------------
//  功能描述 : 针对指令存储器模块 imem 的简单仿真平台
//             • 产生 10 ns 周期、50 % 占空比的 clka
//             • 逐字节地址递增地访问 64 × 32‑bit ROM（0 → 252）
//             • 每次地址变动后立刻打印 rd（验证异步读 / 同步 ROM IP 都兼容）
// ----------------------------------------------------------------------------
//  Verilog‑2001:
//    ‧ 激励 reg，采样 wire。
//    ‧ 主循环写在一个 initial 里，方便扩展为随机地址/特定指令比对。
// ============================================================================

module tb_imem;

  //--------------------------------------------------------------------------
  // DUT 接口
  //--------------------------------------------------------------------------
  reg         clka = 1'b0;  // 仿真主时钟
  reg  [31:0] addr = 32'd0;  // 字节地址输入
  wire [31:0] rd;  // 指令字输出

  //--------------------------------------------------------------------------
  // 被测设计实例化
  //--------------------------------------------------------------------------
  imem dut (
    .clka(clka),
    .a   (addr),
    .rd  (rd)
  );

  //--------------------------------------------------------------------------
  // ① 时钟：10 ns 周期
  //--------------------------------------------------------------------------
  always #5 clka <= ~clka;

  //--------------------------------------------------------------------------
  // ② 主测试流程：线性遍历 ROM 地址
  //--------------------------------------------------------------------------
  integer i;
  initial begin
    // 等待一个正沿，保证 IP 内部逻辑稳定
    @(posedge clka);

    $display("================ IMEM DUMP START ================");

    for (i = 0; i < 64; i = i + 1) begin
      addr <= i;  // 字地址 → 字节地址
      // 等半周期，再取数据（异步 ROM 立即生效；同步 ROM 下一拍生效）
      //#1;  // 1 ns 观察异步效果
      $display("%0t ns : addr = %0h  rd = %0h", $time, addr, rd);
      @(posedge clka);  // 下一拍继续
    end

    $display("================ IMEM DUMP END ==================");
  end

endmodule
