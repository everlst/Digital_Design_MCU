// ============================================================================
//  文件名   : datapath.v
//  模块名   : datapath
//  功能描述 : ARM 单周期 CPU 的 **数据通路**
//             ─ 负责完成指令取址、寄存器读写、立即数扩展、ALU 运算、
//               以及分支 / 跳转目标地址计算。
//             ─ 与 controller 交换控制信号，与外部存储器交换数据。
//             ─ 新增 **Shifter**：支持 Instr[11:5] 所定义的 LSL/LSR/ASR/ROR
//               寄存器移位立即数；结果送 ALU 的 SrcB。
// ----------------------------------------------------------------------------
//  Verilog-2001 迁移要点
//    • 纯组合连线均用 wire；本模块仅例化子模块 + flopr 寄存器。
//    • 端口与旧版保持一致，无接口破坏。
// ----------------------------------------------------------------------------
//  端口列表与说明同旧版，唯独 mux2.d0 由 **WriteData → ShiftedData**。
// ============================================================================
module datapath (
  input clk,
  input reset,

  // ==== 来自 controller 的控制信号 =====================================
  input [1:0] RegSrc,      // 读端口寄存器号来源
  input       RegWrite,    // 寄存器写使能
  input [2:0] ImmSrc,      // 立即数扩展控制
  input       ALUSrc,      // ALU SrcB 选择
  input [2:0] ALUControl,  // ALU 运算控制
  input       MemtoReg,    // 写回数据选择
  input       PCSrc,       // PC 源选择 (顺序 / 跳转)

  // ==== 与 controller 的状态返回 =======================================
  output [3:0] ALUFlags,  // N Z C V

  // ==== 与指令存储器接口 ===============================================
  output [31:0] PC,    // 程序计数器
  input  [31:0] Instr, // 取回的指令

  // ==== 与数据存储器接口 ===============================================
  output [31:0] ALUResult,  // 地址 (STR/LDR) 或运算结果
  output [31:0] WriteData,  // 写入数据存储器的数值 (原始 Rm)
  input  [31:0] ReadData    // 从存储器读出的数据
);

  // --------------------------------------------------------------------
  // 内部连线
  // --------------------------------------------------------------------
  wire [31:0] PCNext, PCPlus4, PCPlus8;  // PC 相关
  wire [31:0] ExtImm;  // 扩展后的立即数
  wire [31:0] SrcA, SrcB;  // 送往 ALU 的两路操作数
  wire [31:0] Result;  // 写回寄存器堆的最终结果
  wire [3:0] RA1, RA2;  // 寄存器堆读端口号
  wire [31:0] ShiftedData;  // Shifter 输出

  // =========================================================================
  // 1) 程序计数器 PC
  // =========================================================================
  mux2 #(
    .WIDTH(32)
  ) pcmux (
    .d0(PCPlus4),
    .d1(Result),
    .s (PCSrc),
    .y (PCNext)
  );

  flopr #(
    .WIDTH(32)
  ) pcreg (
    .clk  (clk),
    .reset(reset),
    .d    (PCNext),
    .q    (PC)
  );

  adder #(
    .WIDTH(32)
  ) pcadd1 (
    .a(PC),
    .b(32'h4),
    .y(PCPlus4)
  );
  adder #(
    .WIDTH(32)
  ) pcadd2 (
    .a(PCPlus4),
    .b(32'h4),
    .y(PCPlus8)
  );

  // =========================================================================
  // 2) 寄存器堆读端口号选择
  // =========================================================================
  mux2 #(
    .WIDTH(4)
  ) ra1mux (
    .d0(Instr[19:16]),
    .d1(4'b1111),
    .s (RegSrc[0]),
    .y (RA1)
  );

  mux2 #(
    .WIDTH(4)
  ) ra2mux (
    .d0(Instr[3:0]),
    .d1(Instr[15:12]),
    .s (RegSrc[1]),
    .y (RA2)
  );

  regfile rf (
    .clk(clk),
    .we3(RegWrite),
    .ra1(RA1),
    .ra2(RA2),
    .wa3(Instr[15:12]),
    .wd3(Result),
    .r15(PCPlus8),
    .rd1(SrcA),
    .rd2(WriteData)      // 未移位的原始 Rm
  );

  // =========================================================================
  // 3) 立即数扩展
  // =========================================================================
  extend ext (
    .Instr (Instr[23:0]),
    .ImmSrc(ImmSrc),
    .ExtImm(ExtImm)
  );

  // =========================================================================
  // 4) **Shifter** ─ 根据 Instr[11:5] 对 WriteData(Rm) 进行移位
  //       shamt = Instr[11:7] (imm5)
  //       shtype = Instr[6:5] (00 LSL / 01 LSR / 10 ASR / 11 ROR)
  // =========================================================================
  shifter shift_u (
    .data_in (WriteData),
    .shamt   (Instr[11:7]),
    .sh_type (Instr[6:5]),
    .data_out(ShiftedData)
  );

  // =========================================================================
  // 5) ALU 第二操作数选择
  //     d0 ← 移位器输出 (寄存器型)
  //     d1 ← 扩展立即数 (立即数型)
  // =========================================================================
  mux2 #(
    .WIDTH(32)
  ) srcbmux (
    .d0(ShiftedData),
    .d1(ExtImm),
    .s (ALUSrc),
    .y (SrcB)
  );

  // =========================================================================
  // 6) ALU
  // =========================================================================
  alu alu_u (
    .a         (SrcA),
    .b         (SrcB),
    .ALUControl(ALUControl),
    .Result    (ALUResult),
    .ALUFlags  (ALUFlags)
  );

  // =========================================================================
  // 7) 写回阶段 MUX
  // =========================================================================
  mux2 #(
    .WIDTH(32)
  ) resmux (
    .d0(ALUResult),
    .d1(ReadData),
    .s (MemtoReg),
    .y (Result)
  );

endmodule
