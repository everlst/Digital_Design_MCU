(* dont_touch = "true" *) module mux3 #(
  parameter WIDTH = 8  // 数据位宽，默认 8 位
) (
  input  [WIDTH-1:0] d0,  // 输入 0
  input  [WIDTH-1:0] d1,  // 输入 1
  input  [WIDTH-1:0] d2,  // 输入 2
  input  [      1:0] s,   // 选择信号（高选 d1，低选 d0）
  output [WIDTH-1:0] y    // 输出
);

  // --------------------------------------------------------------------
  // 组合多路选择：s=0 选 d0，s=1 选 d1
  // --------------------------------------------------------------------


  assign y = (!s[1]) ? (s[0] ? d1 : d0) : d2;

endmodule
