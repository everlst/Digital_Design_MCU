// ============================================================================
//  文件名   : flopenr.v
//  模块名   : flopenr
// ----------------------------------------------------------------------------
//  功能描述 : “带使能、异步复位寄存器”(Flip-Flop with Load-Enable & async Reset)
//             ┌─────────────┐   clk ↑     ┌───────────┐
//             │  输入 d[N:0]├────────────►│           │
//             │  使能 en    │             │   q <= d  │
//             │  复位 reset ├─reset=1───► │   q := 0  │
//             └─────────────┘             └───────────┘
//             • 仅当 en = 1 时才把 d 装载到寄存器；
//             • reset 为高时 **异步** 清零，不受 en 影响；
//             • 位宽由参数 WIDTH 控制，默认 8 位。
// ----------------------------------------------------------------------------
//  Verilog-2001 迁移要点
//    1. SystemVerilog 的 `logic` → Verilog 的 `wire` / `reg`：
//         - q 在时序块内赋值，因此声明为 reg；其余端口默认为 wire。
//    2. 参数列表写法：`#(parameter WIDTH = 8)` **无分号**。
//    3. 时序块用 `always @(posedge clk or posedge reset)` 实现异步复位。
// ============================================================================
module flopenr #(
  parameter WIDTH = 8  // 数据位宽，实例化时可重定义
) (
  input                  clk,    // 时钟
  input                  reset,  // 异步复位（高有效）
  input                  en,     // 载入使能（高采样 d）
  input      [WIDTH-1:0] d,      // 数据输入
  output reg [WIDTH-1:0] q       // 数据输出
);

  // --------------------------------------------------------------------
  // 时序逻辑：异步复位 + 上升沿采样（带使能）
  // --------------------------------------------------------------------
  always @(posedge clk or posedge reset) begin
    if (reset) q <= {WIDTH{1'b0}};  // 复位时立即清零
    else if (en) q <= d;  // 使能为 1 时装载新数据
    // else 保持原值
  end

endmodule
