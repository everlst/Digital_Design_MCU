`timescale 1ns / 1ps
// ============================================================================
//  文件名   : tb_top.v
//  模块名   : tb_top (testbench for top)
// ----------------------------------------------------------------------------
//  功能描述 : 行为级仿真环境，用于验证顶层模块 top
//             ‧ 产生 10 ns 周期、50 % 占空比时钟 clk
//             ‧ 产生同步复位 reset（0 ns–22 ns 高）
//             ‧ 监视 dmem 写端口：
//                • 若向地址 100 写入数据 7  → 输出 **SUCCEEDED** 并结束仿真
//                • 若写地址不是 96（合法的前一次写地址）→ 输出 **FAILED** 并结束仿真
// ----------------------------------------------------------------------------
//  编码规则 : 100 % Verilog‑2001
//             ‧ 激励信号用 reg，DUT 输出用 wire
//             ‧ 所有时序过程赋值使用非阻塞 <=
// ============================================================================

module tb_top;

  //--------------------------------------------------------------------------
  // DUT 接口信号声明
  //--------------------------------------------------------------------------
  reg         clk = 1'b0;  // 系统时钟，0 ns 即确定为 0
  reg         reset;  // 同步复位，高有效
  wire [31:0] WriteData;  // DUT → dmem 写数据
  wire [31:0] DataAdr;  // DUT → dmem 地址
  wire        MemWrite;  // DUT → dmem 写使能

  //--------------------------------------------------------------------------
  // 被测设计实例化
  //--------------------------------------------------------------------------
  top dut (
    .clk  (clk),
    .reset(reset)
    // .WriteData(WriteData),
    // .DataAdr  (DataAdr),
    // .MemWrite (MemWrite)
  );

  //--------------------------------------------------------------------------
  // ① 时钟生成：10 ns 周期，50 % 占空比
  //--------------------------------------------------------------------------
  always #5 clk <= ~clk;

  //--------------------------------------------------------------------------
  // ② 复位脉冲：0 ns–22 ns 为高
  //--------------------------------------------------------------------------
  initial begin
    reset = 1'b1;
    repeat (3) @(posedge clk);  // 至少保持 3 个时钟周期
    reset = 1'b0;  // 退出复位，完全对齐 posedge
  end


  //--------------------------------------------------------------------------
  // ③ 写端口监视与判定逻辑
  //--------------------------------------------------------------------------
  initial begin : WATCH_DMEM_WRITE
    // 等待复位解除再开始监视
    @(negedge reset);

    forever begin
      @(posedge clk);
      if (MemWrite) begin
        $display("%0t ns : Write @ %0d = %0d", $time, DataAdr, WriteData);

        // 成功条件
        if (DataAdr == 32'd100 && WriteData == 32'd7) begin
          $display("\n==================== TEST SUCCEEDED ====================\n");
          // #10 $finish;
        end  // 失败条件
        else if (DataAdr != 32'd96) begin
          $display("\n!!!!!!!!!!!!!!!!!!!! TEST FAILED !!!!!!!!!!!!!!!!!!!!\n");
          // #10 $finish;
        end
        // 其余情况（合法写 96）继续观察
      end
    end
  end


endmodule
