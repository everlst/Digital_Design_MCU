//====================================================================
// 32-bit ALU  (Verilog-2001)
// ────────────────────────────────────────────────────────────────────
// ALUControl[1:0]
//   00 : a + b
//   01 : a - b   (用 ~b + 1 实现二补减法)
//   10 : a & b
//   11 : a | b
// ALUFlags = {N, Z, C, V}
//   N : 结果最高位         (Negative)
//   Z : 结果是否为 0       (Zero)
//   C : 加/减运算产生进位  (Carry)           ─ 仅在加/减时有效
//   V : 加/减运算溢出标志  (Overflow, 2's  complement) ─ 仅在加/减时有效
//====================================================================
module alu (
  input  wire [31:0] a,
  input  wire [31:0] b,
  input  wire [ 1:0] ALUControl,
  output reg  [31:0] Result,      // 用 reg，因为在 always 块里赋值
  output wire [ 3:0] ALUFlags
);

  //----------------------------------------------------------------
  // ① 条件求反 b，再做一条 33-bit 加法得到 sum_ext
  //----------------------------------------------------------------
  wire [31:0] condinvb = (ALUControl[0]) ? ~b : b;  // 01->sub 时取反
  wire [32:0] sum_ext = {1'b0, a} + {1'b0, condinvb} + ALUControl[0];
  wire [31:0] sum = sum_ext[31:0];
  wire        carry_add = sum_ext[32];  // 33-位进位

  //----------------------------------------------------------------
  // ② 根据 ALUControl 产生 Result
  //----------------------------------------------------------------
  always @* begin
    case (ALUControl)
      2'b10:   Result = a & b;
      2'b11:   Result = a | b;
      default: Result = sum;  // 00(add) or 01(sub)
    endcase
  end

  //----------------------------------------------------------------
  // ③ 计算标志位
  //----------------------------------------------------------------
  wire neg = Result[31];  // N
  wire zero = (Result == 32'b0);  // Z
  wire carry = (ALUControl[1] == 1'b0)  // 仅在 add/sub 时有效
  & carry_add;  // C
  wire overflow = (ALUControl[1] == 1'b0)  // 仅在 add/sub 时有效
  & ~(a[31] ^ b[31] ^ ALUControl[0])  // 前两数同号
  & (a[31] ^ Result[31]);  // 与结果异号  → V

  assign ALUFlags = {neg, zero, carry, overflow};
endmodule
