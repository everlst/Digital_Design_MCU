// ==============================================================
//  Arm 5‑Stage Pipeline – Verilog‑2001 Implementation (draft v1)
//  所有模块均保持 Verilog‑2001 语法，已把单周期逻辑改为五级流水，
//  并集成现有 hazard.v（前递+停顿）模块。
//  文件之间用 ----- <filename> ----- 分隔，方便拆分保存。
// ==============================================================

// ------------------------------------------------------------------
// ----- pipeline_top.v --------------------------------------------
// ------------------------------------------------------------------
// SoC 顶层保持不变，只把单周期 CPU 实例替换成 arm_pipeline
// ------------------------------------------------------------------

module pipeline_top (
  input  wire        clk,
  input  wire        rst,
  output wire [31:0] imem_addr,
  input  wire [31:0] imem_rdata,
  output wire [31:0] dmem_addr,
  output wire [31:0] dmem_wdata,
  output wire        dmem_we,
  input  wire [31:0] dmem_rdata
);

  // ---------------------------------------------------------------
  // 实例化五级流水 CPU
  // ---------------------------------------------------------------
  arm_pipeline cpu (
    .clk       (clk),
    .rst       (rst),
    .imem_addr (imem_addr),
    .imem_rdata(imem_rdata),
    .dmem_addr (dmem_addr),
    .dmem_wdata(dmem_wdata),
    .dmem_we   (dmem_we),
    .dmem_rdata(dmem_rdata)
  );

endmodule





// ------------------------------------------------------------------
// ----- hazard.v (保持接口一致，内部逻辑已在原文件) --------------
// ------------------------------------------------------------------
// 如需调整可在此文件修改；本示例假设原 hazard.v 逻辑符合接口

// ------------------------------------------------------------------
// 其余模块 (alu.v, extend.v, regfile.v, adder.v, mux2.v, flopr.v 等)
// 均保持原单周期版本，可直接复用。
// ------------------------------------------------------------------

// ==============================================================
//  End of File
// ==============================================================
