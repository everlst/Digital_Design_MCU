// ============================================================================
//  文件名   : extend.v
//  模块名   : extend
// -----------------------------------------------------------------------------
//  功能描述 : 立即数扩展单元（ARM 单周期 CPU）
//             ─ 根据控制信号 ImmSrc[1:0] 选择不同的扩展方式，
//               生成 32-bit 立即数 ExtImm 送往 ALU / 地址计算。
// -----------------------------------------------------------------------------
//  Verilog-2001 版本说明
//    • SystemVerilog 的  logic / always_comb → Verilog 的 reg / always @*。
//    • 输出 ExtImm 在组合 always 块内赋值，故声明为 reg 类型。
// -----------------------------------------------------------------------------
(* dont_touch = "true" *) module extend (
  input      [23:0] Instr,   // 指令位段 (不同指令使用位宽不同的立即数字段)
  input      [ 2:0] ImmSrc,  // 立即数来源选择
  output reg [31:0] ExtImm   // 扩展后的 32-bit 立即数
);

  // =========================================================================
  // 立即数扩展规则
  // -------------------------------------------------------------------------
  // ImmSrc = 00 : 数据处理指令  —— 取 Instr[7:0]，零扩展到 32 位
  // ImmSrc = 01 : LDR/STR 偏移  —— 取 Instr[11:0]，零扩展到 32 位
  // ImmSrc = 10 : Branch 偏移   —— 取 Instr[23:0]，先带符号扩展到 28 位，
  //                                再左移 2 位补 2 个零，形成 32 位偏移
  // 其它值       : 未定义，输出 X
  // =========================================================================
 (* dont_touch = "true" *) wire [4:0] sh = {Instr[11:8], 1'b0};  // rot*2
 (* dont_touch = "true" *)  reg  [7:0] Temp;

  always @* begin
    case (ImmSrc)
      3'b000:  ExtImm = {24'b0, Instr[7:0]};  // 8 位零扩展
      3'b001:  ExtImm = {20'b0, Instr[11:0]};  // 12 位零扩展
      3'b010:  ExtImm = {{6{Instr[23]}}, Instr[23:0], 2'b00};  // 24 位有符号扩展再左移 2
      3'b011: begin
        Temp   = {Instr[7:0], Instr[7:0]} >> sh;
        ExtImm = {24'b0, Temp[7:0]};
      end
      default: ExtImm = 32'bx;  // 未定义
    endcase
  end

endmodule
