// ============================================================================
//  文件名   : flopr.v
//  模块名   : flopr
// ----------------------------------------------------------------------------
//  功能描述 : “同步复位寄存器”（Flip-Flop with synchronous Reset）
//             ─ 宽度可参数化，默认 8 位。
//             ─ 在时钟上升沿采样 d；若 reset=1，则输出 q 被清零。
//             ─ 常用于流水线寄存器、程序计数器等需要同步复位的场合。
// ----------------------------------------------------------------------------
//  Verilog-2001 编码要点
//    1. SystemVerilog 的 `logic` → Verilog 的 `reg` / `wire`。
//       · 本例中 q 在时序块内赋值，声明为 reg。
//       · clk、reset、d 仅作输入连线，省略类型默认为 wire。
//    2. `always_ff` 换成传统时序块 `always @(posedge clk)`；
//       同步复位需在时序内用 if…else 判断。
//    3. ANSI-style 端口写法（IEEE-1364-2001）已经支持大多数工具链。
// ----------------------------------------------------------------------------
(*DONT_TOUCH="YES"*) module flopr #(
  parameter WIDTH = 8  // 数据位宽（可在实例化时重定义）
) (
  input                  clk,    // 时钟
  input                  reset,  // 同步复位（高有效）
  input      [WIDTH-1:0] d,      // 数据输入
  output reg [WIDTH-1:0] q       // 数据输出
);

  // --------------------------------------------------------------------
  // 时序逻辑：同步复位 + 边沿采样
  // --------------------------------------------------------------------
  always @(posedge clk or posedge reset) begin
    if (reset) q <= 0;  // 复位时清零
    else q <= d;  // 采样输入
  end

endmodule
