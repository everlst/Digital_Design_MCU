// ============================================================================
//  文件名   : adder.v
//  模块名   : adder
// ----------------------------------------------------------------------------
//  功能描述 : 可参数化位宽的纯组合加法器
//             ┌────────────┐      ┌────────────┐
//             │ 输入 a[N:0]│ ---> │            │
//             │ 输入 b[N:0]│ ---> │   y = a+b  │ ---> 输出 y[N:0]
//             └────────────┘      └────────────┘
//             • 结果 y 与输入位宽相同，若溢出则高位被截断。
//             • 完全组合逻辑（assign），综合后映射为加法器或查找表。
// ----------------------------------------------------------------------------
//  Verilog-2001 说明
//    1. SystemVerilog 写法 `parameter WIDTH = 8;` 末尾分号需删除：
//         → `#(parameter WIDTH = 8)`
//    2. 去除 `logic` 关键字，端口未显式声明类型时默认为 wire。
//    3. `always_comb` 替换为连续赋值 `assign`，避免使用 reg。
// ============================================================================
 module adder #(
  parameter WIDTH = 8  // 数据位宽，默认 8 位
) (
  input  [WIDTH-1:0] a,  // 加数
  input  [WIDTH-1:0] b,  // 被加数
  output [WIDTH-1:0] y   // 求和结果
);

  // --------------------------------------------------------------------
  // 纯组合加法：工具会综合为硬件加法器或 LUT
  // --------------------------------------------------------------------
  assign y = a + b;

endmodule
