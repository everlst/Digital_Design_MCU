// ==============================================================
//  Arm 5-Stage Pipeline – Verilog-2001 Implementation (draft v2)
//  更新内容：
//    • 新增 SoC 顶层  soc_top.v   —— 连接 ROM(IP) + dmem + arm_pipeline
//    • 行为级 ROM (imem_rom.v)   —— 如不用，可替换成厂商 Block‑ROM IP
//    • 简易 TestBench  tb_soc.v  —— 时钟、复位、VCD 波形、运行 5 µs
//  其余文件（arm_pipeline.v、controller.v、hazard.v…）沿用 v1 版本
// ==============================================================

// ------------------------------------------------------------------
// ----- soc_top.v ---------------------------------------------------
// ------------------------------------------------------------------
// 顶层：ROM → 指令流， dmem → 数据流， CPU = arm_pipeline
// ------------------------------------------------------------------
module soc_top (
  input wire clk,
  input wire rst
);

  // ---------------- CPU ↔ 指令存储器 -----------------------------
  wire [31:0] imem_addr;
  wire [31:0] imem_rdata;

  // ---------------- CPU ↔ 数据存储器 -----------------------------
  wire [31:0] dmem_addr;
  wire [31:0] dmem_wdata;
  wire        dmem_we;
  wire [31:0] dmem_rdata;

  // ---------------------------------------------------------------
  // 行为级指令 ROM（如用 Xilinx/Intel IP，可直接实例化 IP 核）
  // ---------------------------------------------------------------
  // 指令存储器（仿真只读 ROM）
  //    • 读延迟 0，地址直接为 PC（字地址对齐）  
  //    • 端口惯例：.a → address, .rd → read-data
  // =========================================================================
  imem im (
    .clka(clk),        // 时钟
    .a   (imem_addr),
    .rd  (imem_rdata)
  );

  // ---------------------------------------------------------------
  // 数据存储器：延用原 dmem.v（双口 RAM/单口 RAM 均可）
  // ---------------------------------------------------------------
  dmem u_dmem (
    .clk(clk),
    .we (dmem_we),
    .a  (dmem_addr),
    .wd (dmem_wdata),
    .rd (dmem_rdata)
  );

  // ---------------------------------------------------------------
  // 5‑级流水 CPU
  // ---------------------------------------------------------------
  arm_pipeline cpu (
    .clk       (clk),
    .rst       (rst),
    .imem_addr (imem_addr),
    .imem_rdata(imem_rdata),
    .dmem_addr (dmem_addr),
    .dmem_wdata(dmem_wdata),
    .dmem_we   (dmem_we),
    .dmem_rdata(dmem_rdata)
  );

endmodule
