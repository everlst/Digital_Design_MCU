// ============================================================================
//  文件名   : dmem.v
//  模块名   : dmem
// ----------------------------------------------------------------------------
//  功能描述 : **32-bit 单端口数据存储器**（写同步、读异步）  
//             • 地址宽度 64 × 4 Byte  → 256 Byte（可按需扩展）  
//             • 地址 a[31:2] 作为字地址（低 2 位舍弃，统一字对齐）  
//             • 写操作：posedge clk 时，若 we=1 把 wd 写入 RAM[…]  
//             • 读操作：异步组合，rd = RAM[…]                   │
// ----------------------------------------------------------------------------
//  Verilog-2001 迁移要点
//    1. SystemVerilog 的 `logic` → Verilog 的 `reg` / `wire`  
//       · 内部阵列 `RAM`、输出 `rd` 在 always 块或 assign 中赋值，需 `reg`。  
//    2. `always_ff` → `always @(posedge clk)`（同步写）  
//    3. ANSI-style 端口使用 IEEE-1364-2001 语法，综合工具普遍支持。  
// ============================================================================
module dmem (
  input         clk,  // 时钟
  input         we,   // 写使能（高有效）
  input  [31:0] a,    // 地址（字节对齐，取高位[31:2] 作索引）
  input  [31:0] wd,   // 写入数据
  output [31:0] rd    // 读出数据
);

  // --------------------------------------------------------------------
  // 1) 内部存储阵列：64 × 32-bit（可通过修改深度扩展容量）
  // --------------------------------------------------------------------
  // reg [31:0] RAM[63:0];  // RAM[0]…RAM[63] ↔ 地址范围 0x00–0xFC
  reg [15:0] RAM[256:0];
  // 行为级仿真初始化
  initial begin
    // ① 如果你已经有一个纯 HEX / BIN 列表：
    $readmemh("FFT_input.mem", RAM);  // 每行一字（16-bit）
  end

  // --------------------------------------------------------------------
  // 2) 异步读：地址变化即刻输出
  // --------------------------------------------------------------------

  // assign rd = RAM[a[31:2]];  // 舍弃最低 2 位，实现字对齐
  assign rd = RAM[a[8:1]];

  // --------------------------------------------------------------------
  // 3) 同步写：上升沿写入
  // --------------------------------------------------------------------
  always @(posedge clk) begin
    // if (we) RAM[a[31:2]] <= wd;
    if (we) RAM[a[8:1]] <= wd;
  end

endmodule
