// ============================================================================
//  文件名   : regfile.v
//  模块名   : regfile
// -----------------------------------------------------------------------------
//  功能描述 : 16 × 32-bit 通用寄存器堆（单写双读）
///           • R0  ─ R14 存放于片上寄存器阵列 rf[0:14]                      │
///           • R15 (PC) 由外部连线 r15 提供，不写入阵列                    │
///           • 每个时钟上升沿，若 we3=1 则把 wd3 写入 wa3 所指定的寄存器    │
///           • 两个读端口 ra1 / ra2 为组合输出；若索引=15 则直接返回 r15   │
// -----------------------------------------------------------------------------
//  Verilog-2001 注意事项
//    1. SystemVerilog 的 `logic` / `always_ff` 改为 Verilog `reg` / `always`
//    2. `reg [31:0] rf [0:14];` 的数组索引从 0—14，对应 R0–R14
//    3. 输出端口 rd1/rd2 在连续赋值下默认为 wire 类型（无须额外声明）
// ============================================================================
 module regfile (
  input         clk,  // 时钟
  input         we3,  // 写使能（高有效）
  input  [ 3:0] ra1,  // 读端口 A 寄存器号
  input  [ 3:0] ra2,  // 读端口 B 寄存器号
  input  [ 3:0] wa3,  // 写端口寄存器号
  input  [31:0] wd3,  // 写入数据
  input  [31:0] r15,  // 外部提供的 PC 值 (R15)
  output [31:0] rd1,  // 读端口 A 数据
  output [31:0] rd2   // 读端口 B 数据
);

  // --------------------------------------------------------------------
  // 16 × 32-bit 寄存器阵列（仅存储 R0–R14，共 15 个槽位）
  // --------------------------------------------------------------------
   reg [31:0] rf[14:0];  // rf[0]↔R0 … rf[14]↔R14

  // --------------------------------------------------------------------
  // 同步写端口
  //   • 每逢 clk 上升沿，若 we3=1 /////////////////////////////////////////////////////且 wa3≠15，则更新对应寄存器
  //   • 若 wa3 为 15（PC），按 ARM 规范应由外部逻辑处理；此处忽略写
  // --------------------------------------------------------------------
  always @(posedge clk) begin
    if (we3 && wa3 != 4'd15)  // 加一条写保护
      rf[wa3] <= wd3;
  end


  // --------------------------------------------------------------------
  // 组合读端口
  //   • 如果索引 = 15 则直接返回 r15 (PC+8)                    │
  //   • 否则从阵列中取值                                     │
  // --------------------------------------------------------------------
  assign rd1 = (ra1 == 4'b1111) ? r15 : rf[ra1];  // 读端口 A
  assign rd2 = (ra2 == 4'b1111) ? r15 : rf[ra2];  // 读端口 B

endmodule
